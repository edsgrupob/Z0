-- Elementos de Sistemas
-- by Luciano Soares
-- Register8.vhd

Library ieee; 
use ieee.std_logic_1164.all;
  
entity Register8 is
	port(
		clock:   in STD_LOGIC;
		input:   in STD_LOGIC_VECTOR(7 downto 0);
		load:    in STD_LOGIC;
		output: out STD_LOGIC_VECTOR(7 downto 0)
	);
end entity;

architecture arch_Register8 of Register8 is

component BinaryDigit
	port(
		clock:   in STD_LOGIC;
		input:   in STD_LOGIC;
		load:    in STD_LOGIC;
		output: out STD_LOGIC
	);
end component;

begin 
	u1: BinaryDigit port map (clock, input, load, output);
	u2: BinaryDigit port map (clock, input, load, output);
	u3: BinaryDigit port map (clock, input, load, output);
	u4: BinaryDigit port map (clock, input, load, output);
	u5: BinaryDigit port map (clock, input, load, output);
	u6: BinaryDigit port map (clock, input, load, output);
	u7: BinaryDigit port map (clock, input, load, output);
	u8: BinaryDigit port map (clock, input, load, output);
end architecture;